(** printing |-#    %\vdash_{\#}%    #&vdash;<sub>&#35;</sub>#     *)
(** printing |-##   %\vdash_{\#\#}%  #&vdash;<sub>&#35&#35</sub>#  *)
(** printing |-##v  %\vdash_{\#\#v}% #&vdash;<sub>&#35&#35v</sub># *)
(** printing |-!    %\vdash_!%       #&vdash;<sub>!</sub>#         *)
(** remove printing ~ *)

Set Implicit Arguments.

Require Import LibLN.
Require Import Coq.Program.Equality.
Require Import Definitions.
Require Import Narrowing.
Require Import Helper_lemmas.
Require Import Precise_types.

(** This module contains lemmas related to invertible typing
    ([ty_var_inv], [|-##] and [ty_val_inv], [|-##v]). *)

(** Invertible-to-precise typing for field declarations: #<br>#
    [Gamma |-## x: {a: T}]
    ----------------------
    [exists T'. Gamma |-! x: {a: T'}]      #<br>#
    [Gamma |-# T' <: T]. *)
Lemma invertible_to_precise_trm_dec: forall G x a T,
  G |-## x : typ_rcd (dec_trm a T) ->
  exists T',
    G |-! trm_var (avar_f x) : typ_rcd (dec_trm a T') /\
    G |-# T' <: T.
Proof.
  introv Hinv.
  dependent induction Hinv.
  - exists T. auto.
  - specialize (IHHinv _ _ eq_refl). destruct IHHinv as [V [Hx Hs]].
    exists V. split; auto.
    eapply subtyp_trans_t; eassumption.
Qed.

(** Invertible-to-precise typing for function types: #<br>#
    [ok Gamma]                        #<br>#
    [Gamma |-## x: forall(S)T]
    ----------------------
    [exists S', T'. Gamma |-! x: forall(S')T']  #<br>#
    [Gamma |-# S <: S']               #<br>#
    [Gamma |-# T'^y <: T^y], where [y] is fresh. *)
Lemma invertible_to_precise_typ_all: forall G x S T,
  ok G ->
  G |-## x : typ_all S T ->
  exists S' T' L,
    G |-! trm_var (avar_f x) : typ_all S' T' /\
    G |-# S <: S' /\
    (forall y,
        y \notin L ->
            G & y ~ S |- open_typ y T' <: open_typ y T).
Proof.
  introv HG Hinv.
  dependent induction Hinv.
  - exists S T (dom G); auto.
  - specialize (IHHinv _ _ HG eq_refl).
    destruct IHHinv as [S' [T' [L' [Hpt [HSsub HTsub]]]]].
    exists S' T' (dom G \u L \u L').
    split; auto.
    assert (Hsub2 : G |-# typ_all S0 T0 <: typ_all S T).
    { apply subtyp_all_t with (L:=L); assumption. }
    split.
    + eapply subtyp_trans_t; eauto.
    + intros y Fr.
      assert (Hok: ok (G & y ~ S)) by auto using ok_push.
      apply tight_to_general in H; auto.
      assert (Hnarrow: G & y ~ S |- open_typ y T' <: open_typ y T0).
      { eapply narrow_subtyping; auto using subenv_last. }
      eauto.
Qed.

(** * Invertible Variable Typing *)

(** Invertible typing is closed under tight subtyping. *)
Lemma invertible_typing_closure_tight: forall G x T U,
  inert G ->
  G |-## x : T ->
  G |-# T <: U ->
  G |-## x : U.
Proof.
  intros G x T U Hgd HT Hsub.
  dependent induction Hsub; eauto.
  - inversion HT.
    destruct (precise_bot_false Hgd H).
  - inversion HT; auto. apply ty_and1_p in H. auto.
  - inversion HT; auto. apply ty_and2_p in H. auto.
  - inversions HT.
    + false* precise_psel_false.
    + pose proof (inert_unique_tight_bounds Hgd H H5) as Hu. subst. assumption.
Qed.

(** ** Tight-to-Invertible Lemma for Variables

       This lemma corresponds to Theorem 3.6 in the paper.

       [inert Gamma]            #<br>#
       [Gamma |-# x: U]
       -----------------
       [Gamma |-## x: U] *)
Lemma tight_to_invertible :
  forall G U x,
    inert G ->
    G |-# trm_var (avar_f x) : U ->
    G |-## x : U.
Proof.
  intros G U x Hgd Hty.
  dependent induction Hty.
  - auto.
  - specialize (IHHty _ Hgd eq_refl).
    eapply ty_bnd_inv.
    apply IHHty.
  - specialize (IHHty _ Hgd eq_refl).
    inversion IHHty; subst; auto.
  - apply ty_and_inv; auto.
  - eapply invertible_typing_closure_tight; auto.
Qed.

(** * Invertible Value Typing *)

(** Invertible value typing is closed under tight subtyping. *)
Lemma invertible_typing_closure_tight_v: forall G v T U,
  inert G ->
  G |-##v v : T ->
  G |-# T <: U ->
  G |-##v v : U.
Proof.
  introv Hgd HT Hsub.
  dependent induction Hsub; eauto; inversions HT; auto; try solve [inversion* H].
  - inversions H0.
  - lets Hb: (inert_unique_tight_bounds Hgd H H5). subst*.
Qed.

(** ** Tight-to-Invertible Lemma for Values

       [inert Gamma]            #<br>#
       [Gamma |-# v: T]
       -----------------
       [Gamma |-##v v: T] *)
Lemma tight_to_invertible_v : forall G v T,
    inert G ->
    G |-# trm_val v : T ->
    G |-##v v : T.
Proof.
  introv Hgd Hty.
  dependent induction Hty; eauto.
  specialize (IHHty v Hgd eq_refl).
  apply* invertible_typing_closure_tight_v.
Qed.
